library verilog;
use verilog.vl_types.all;
entity ula_32bit_vlg_vec_tst is
end ula_32bit_vlg_vec_tst;
