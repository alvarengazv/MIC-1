library verilog;
use verilog.vl_types.all;
entity DATA_PATH_vlg_vec_tst is
end DATA_PATH_vlg_vec_tst;
