library verilog;
use verilog.vl_types.all;
entity MAR is
    port(
        DATA_ADDRESS    : out    vl_logic_vector(31 downto 0);
        LOAD            : in     vl_logic;
        MIR             : in     vl_logic_vector(35 downto 0);
        CLOCK           : in     vl_logic;
        IN_C            : in     vl_logic_vector(31 downto 0)
    );
end MAR;
