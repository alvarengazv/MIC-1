library verilog;
use verilog.vl_types.all;
entity MBR_EXTENSOR_vlg_vec_tst is
end MBR_EXTENSOR_vlg_vec_tst;
